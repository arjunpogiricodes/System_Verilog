


// class inheritance and constrint overidden
// grandparent class declaration

class grandparent;
         randc int pkt1;
         constraint over_pkt1{ pkt1 > 50;}
         randc int pkt2;
         constraint over_pkt2{ pkt2 < 50 ;}
         randc int  pkt3;
         constraint over_pkt3{ pkt3 > 50 && pkt3 < 200;}
         randc int pkt4;
         constraint over_pkt4{ pkt4 > 50 && pkt4 < 150;}

         function void  post_randomize;
               $display("\n***************************** grand parent class *********************************************\n");
               $display("pkt1 = %0d type = %s \npkt2 = %0d  type = %s \npkt3 = %0d type = %s \npkt4 = %0d type = %s",pkt1,$typename(pkt1),pkt2,$typename(pkt2),pkt3,$typename(pkt3),pkt4,$typename(pkt4));
               $display("\n******************************************************************************************\n");
         endfunction:post_randomize 

     
endclass:grandparent

// parent class  declaration

class parent extends grandparent;
            
         //bit[7:0] pkt1;
         constraint under_pkt1{ pkt1 < 150;}
         //rand bit[7:0] pkt2;
         constraint over_pkt2{ (pkt2  > 50) && (pkt2 < 150);}
         randc bit[7:0] pkt3;
         constraint over_pkt3{ pkt3  < 50;}
         randc bit[7:0] pkt4;
         constraint under_pkt4{ pkt4 > 100;}

         function void  post_randomize;
               $display("\n***************************** parent class *********************************************\n");
               $display("pkt1 = %0d type = %s \npkt2 = %0d  type = %s \npkt3 = %0d type = %s \npkt4 = %0d type = %s",pkt1,$typename(pkt1),pkt2,$typename(pkt2),pkt3,$typename(pkt3),pkt4,$typename(pkt4));
               $display("\n******************************************************************************************\n");
         endfunction:post_randomize 
endclass:parent

// declaring the handles
 
        grandparent ga; 
        parent pa;
       
//creating mdoule

module test;
        
        initial begin 
        ga = new;
        pa = new;
        for(int i= 0;i<10;i++)
           begin
           //ga.randomize;
           pa.randomize; 
           $display("\n#####################################################################################\n");
           $display(" %0p " ,pa);
           $display("\n#####################################################################################\n");
           end
        end

endmodule:test

/*
***************************** parent class *********************************************

pkt1 = 98 type = int 
pkt2 = 126  type = int 
pkt3 = 25 type = bit[7:0] 
pkt4 = 124 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:98, pkt2:126, pkt3:-1559125241, pkt4:66, pkt3:'h19, pkt4:'h7c} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 147 type = int 
pkt2 = 117  type = int 
pkt3 = 8 type = bit[7:0] 
pkt4 = 142 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:147, pkt2:117, pkt3:1369010820, pkt4:149, pkt3:'h8, pkt4:'h8e} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 91 type = int 
pkt2 = 64  type = int 
pkt3 = 37 type = bit[7:0] 
pkt4 = 239 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:91, pkt2:64, pkt3:2035665862, pkt4:134, pkt3:'h25, pkt4:'hef} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 58 type = int 
pkt2 = 77  type = int 
pkt3 = 45 type = bit[7:0] 
pkt4 = 211 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:58, pkt2:77, pkt3:1832097639, pkt4:52, pkt3:'h2d, pkt4:'hd3} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 102 type = int 
pkt2 = 57  type = int 
pkt3 = 19 type = bit[7:0] 
pkt4 = 147 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:102, pkt2:57, pkt3:-1006585545, pkt4:54, pkt3:'h13, pkt4:'h93} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 137 type = int 
pkt2 = 58  type = int 
pkt3 = 42 type = bit[7:0] 
pkt4 = 136 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:137, pkt2:58, pkt3:-1869009377, pkt4:113, pkt3:'h2a, pkt4:'h88} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 90 type = int 
pkt2 = 80  type = int 
pkt3 = 21 type = bit[7:0] 
pkt4 = 207 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:90, pkt2:80, pkt3:-1160387189, pkt4:91, pkt3:'h15, pkt4:'hcf} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 127 type = int 
pkt2 = 81  type = int 
pkt3 = 12 type = bit[7:0] 
pkt4 = 165 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:127, pkt2:81, pkt3:-1342996415, pkt4:76, pkt3:'hc, pkt4:'ha5} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 78 type = int 
pkt2 = 91  type = int 
pkt3 = 33 type = bit[7:0] 
pkt4 = 223 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:78, pkt2:91, pkt3:-1520389468, pkt4:140, pkt3:'h21, pkt4:'hdf} 

#####################################################################################


***************************** parent class *********************************************

pkt1 = 57 type = int 
pkt2 = 133  type = int 
pkt3 = 4 type = bit[7:0] 
pkt4 = 169 type = bit[7:0]

******************************************************************************************


#####################################################################################

 '{pkt1:57, pkt2:133, pkt3:53029846, pkt4:116, pkt3:'h4, pkt4:'ha9} 

#####################################################################################

*/


