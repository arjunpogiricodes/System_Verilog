


// creating interface
// mod 12 up down mode counter

//`define int no_of_gen = 50;

interface inter(input bit clk);

     logic[3:0] data_out;

     bit mode;

     bit reset;

     bit load;

     logic[3:0] data_in;

// cloking block for write driver

   clocking wd_cb@(posedge clk);
        default  input#1 output #1;

           output mode;
           output reset;
	   output load;
	   output data_in;
		  
    endclocking:wd_cb

// clocking block for write monitor

     clocking wm_cb@(posedge clk);
           default input #1 output #1;

             input mode;
             input reset;
	     input load;
	     input data_in;
			 
     endclocking:wm_cb

// clocking block for read monitor 

    clocking rm_cb@(posedge clk);
          default input #1 output #1;

             input mode;
	     input load;
             input data_out;  
             input reset;
			 
     endclocking:rm_cb

     modport WD(clocking wd_cb);
     modport WM(clocking wm_cb);
     modport RM(clocking rm_cb);
     //modport DUV(input clk,input mode,input reset,input load,input data_in,output data_out);

endinterface:inter

module counter(clk,reset,load,mode,data_in,data_out);
 
        input bit clk,mode,reset,load;
        input logic[3:0] data_in;
        output logic[3:0] data_out;
           
    
     always@(posedge clk)
        begin
          
          if(reset == 1'b0)
		  
              data_out <= 4'd0;
			   
          else if(load == 1'b1)
		  
              data_out <= data_in;
				 
          else if(mode == 1'b0)
		  
                if(data_out == 4'd0)
                     data_out <= 4'd11;
                else
                     data_out <= data_out - 1'b1; 
					 
          else if(mode == 1'b1)
		  
               if(data_out >= 4'd11)
                     data_out <= 4'd0;
               else
                     data_out <= data_out +1'b1; 
       end
endmodule:counter

// class trasaction 
class packet;

     logic[3:0] data_out;

      rand bit mode;

      rand bit reset;

      rand bit load ;

      rand logic[3:0] data_in;

          constraint val_data  { data_in inside{[0:11]};}
	  constraint reset_con { reset   dist{ 1'b0:=30,1'b1:=50};}
	  constraint mode_con  { mode    dist{ 1'b0:=20,1'b1:=50};}
	  constraint load_con  { load    dist{ 1'b0:=50,1'b1:=20};}
	  
	  
	  
	  static int no_trans_id;
	  static int no_load;
	  static int no_reset;
	  static int no_mode;
	 

     function void post_randomize();
          
         if(load == 1'b1);
             no_load++;
         if(mode == 1'b1);
             no_mode++;
         if(reset == 1'b0);
             no_reset++;

	 $display("no_load = %0d no_mode = %0d no_reset = %0d ",no_load,no_mode,no_reset);	 
         $display("\n==================================== post randomize  t=%0t ==================================================\n",$time);   
         $display("\n reset = %b load = %b data_in = %0d mode = %b\n",reset,load,data_in,mode); 
         $display("\n==============================================================================================================\n");
      
     endfunction:post_randomize

endclass:packet     

// class generator 

class generator;

        int no_of_gen = 200;
        packet pa,pb;

        mailbox #(packet) ma;

        function new(mailbox #(packet) ma);
               
             this.ma = ma;
              pa = new;
        endfunction:new

        task start();
            for(int i=0; i< no_of_gen;i++)
              begin
                  //pa = new;
				  pa.no_trans_id++;
                  assert(pa.randomize())
                     else $display("\n!!!!!!!!!!!!!!!!!!!!!!!!!!Randomize Violation!!!!!!!!!!!!!!!!!!!!!!!!!!!!\n");
                  pb = new pa;
                  ma.put(pb);
	          $display("\n====================================== generator no_trans_id = %0d======================================\n ",pa.no_trans_id,$time);
              end
        endtask:start

 endclass:generator



class write_drive;

         packet pa,pb;
         virtual inter.WD  wd_inter;
         mailbox #(packet) ma;
		 function new(virtual inter.WD  wd_inter,mailbox #(packet) ma);
		         this.wd_inter = wd_inter;
		         this.ma = ma;
		 endfunction:new
        
		 virtual task drive();
		 
               @(wd_inter.wd_cb);
	       wd_inter.wd_cb.reset   <= pb.reset;
	       wd_inter.wd_cb.mode    <= pb.mode;
	       wd_inter.wd_cb.load    <= pb.load;
	       wd_inter.wd_cb.data_in <= pb.data_in;
             		   
		 endtask:drive
		
         task start();
                fork begin 
                          forever begin
                                ma.get(pa);
				pb = new pa;
                                drive();
			        $display("\n====================================== Write Driver t=%0t ======================================\n ",$time);
                              end
                      end
                join_none
         endtask:start

         		 
endclass:write_drive


// class write monitor

class write_monitor;

          virtual inter.WM wm_inter;
             
          mailbox #(packet) ma;
          packet pa,pb;
           
          function new(	virtual inter.WM wm_inter,mailbox #(packet) ma);
                
                      this.wm_inter = wm_inter;
                      this.ma = ma;
		      pa = new;
					  
          endfunction:new
		  
		   
		  virtual task monitor();

                                 @(wm_inter.wm_cb);
				   begin
				     pa.reset = wm_inter.wm_cb.reset;
				     pa.mode = wm_inter.wm_cb.mode;
				     pa.load = wm_inter.wm_cb.load;
				     pa.data_in = wm_inter.wm_cb.data_in;
				   end
          endtask:monitor
		  
          task start();
		  
		         fork begin
				  forever
				     begin
					 monitor();
				         pb = new pa;
		                         ma.put(pb);
				         $display("\n====================================== Write Monitor t=%0t ======================================\n ",$time);
				          $display(" Reset = %b Mode = %b  Load = %b Data_in  = %0d ",pa.reset,pa.mode,pa.load,pa.data_in);
				         $display("\n=========================================================================================================\n");

          		              end
				    end
		            join_none	   
           endtask:start

endclass:write_monitor


// class read monitor

class read_monitor;

            virtual inter.RM rm_inter;
            mailbox #(packet) ma;
			packet pa,pb;
			
			function new(virtual inter.RM rm_inter,mailbox #(packet) ma);
			
			         this.rm_inter = rm_inter;
					 this.ma = ma;
					 this.pa = new;
		    endfunction:new

            virtual task monitor();
			        @(rm_inter.rm_cb);
			         begin
					 
			         pa.data_out = rm_inter.rm_cb.data_out;
                                 pa.reset = rm_inter.rm_cb.reset; 
                                 pa.load = rm_inter.rm_cb.load; 
                                 pa.mode = rm_inter.rm_cb.mode; 
					 
			         end

             endtask:monitor

            task start();
                  fork begin 
                            forever begin
                                      monitor(); 
				      pb = new pa;
                                      ma.put(pb);
				      $display("\n====================================== Read Monitor t=%0t ======================================\n ",$time);
				      $display(" Reset = %b Mode = %b  Load = %b Data_out  = %0d ",pb.reset,pb.mode,pb.load,pb.data_out);
				      $display("\n=========================================================================================================\n");
                                   end									  
			    end
		   join_none	   
	    endtask:start
			 
endclass:read_monitor

class refence_model;

          packet pa,pb;
          mailbox #(packet) mw,sbm;
	  bit [3:0] data_out;
	  function new(mailbox #(packet) mw,mailbox #(packet) sbm);

	         this.mw = mw;
                 this.sbm = sbm;
				 
	 endfunction:new
	 
	 task model(packet pb);   
        
		if(pb.reset == 1'b0)
		
                     data_out <= 4'd0;
          
		else if(pb.load == 1'b1)
          
        	      data_out <= pb.data_in;
					 
               //wait (pb.load == 1'b0) 
		// begin
 	        else if(pb.mode == 1'b1)           
         
        		if(data_out >= 4'd11)
				
                            data_out <= 4'd0;
					 
                         else
                            data_out <= data_out + 1'b1;  
           
   	        else if(pb.mode == 1'b0)
           
     		       if(data_out == 4'd0)
             
           			 data_out <= 4'd11;
                       else
          
             		 data_out <= data_out - 1'b1;
		 			  
	  
					 
      endtask:model
      	
	  task start();
           fork begin
                     forever
                            begin
			       mw.get(pa);
			       pb = new pa;
			       model(pb);
			       pb.data_out = data_out; 
			     sbm.put(pb);
			     $display("\n====================================== Refence Model t=%0t ======================================\n ",$time);
			     $display(" Reset = %b Mode = %b  Load = %b Data_out  = %0d ",pb.reset,pb.mode,pb.load,pb.data_out);
			     $display("\n=========================================================================================================\n");
								 
			   end 		 

                  end
           join_none
       endtask:start

endclass:refence_model


// score board

class score_board;

        packet prf,prm;
		mailbox #(packet) mrf,mrm;
		string dff;
		int no_compare;
		 event DONE;
		
		function new(mailbox #(packet) mrf,mailbox #(packet) mrm);
		         
				  this.mrf = mrf;
				  this.mrm = mrm;
                                  this.cg = new;       
		endfunction:new

           function void compare(packet prf,packet prm,output string dff);
   			    no_compare++;
                                 cg.sample; 

				if(prf.data_out == prm.data_out ) 
				    begin
                                        
			                dff = "\n##########################################################################################\n\t\t Success Fully Compare \n##########################################################################################\n";
					   //return 1'b1; 
			            end
			         else 
				      begin
                                       dff = "\n##########################################################################################\n\t\t Compare is Failed \n##########################################################################################\n";
                        //return 1'b1; 					
                                       end                    					  
             endfunction:compare

             covergroup  cg;

                     DATA_OUT: coverpoint prm.data_out{
                                                      bins  val1 = {[0:1]};
                                                      bins  val2 = {[2:3]};
                                                      bins  val3 = {[4:5]};
                                                      bins  val4 = {[6:7]};
                                                      bins  val5 = {[7:8]};
                                                      bins  val6 = {[8:9]};
                                                      bins  val7 = {[9:11]};

                                                      }
                     MODE: coverpoint prm.mode{ 
                                                    bins val8[] = {0,1};
                                              }
                     LOAD:  coverpoint prm.load{
                                                      bins val9[] = {0,1};
                                              }
                     RESET: coverpoint prm.reset{
                                                     bins val10[] = {0,1};
                                               } 
                     RXLXMXDO	: cross DATA_OUT,MODE,LOAD;
                     
 
	    endgroup:cg	
 
	     task start();
		    fork begin
			       forever begin
				          mrf.get(prf);
			                  mrm.get(prm);
				          compare(prf,prm,dff);
					  $display(dff);
                                          $display("...............   %f  ................",cg.get_coverage());
                                          if(no_compare == prm.no_trans_id)
					      begin
						 -> DONE;
					       end	
					end
                  end
              join_none
        endtask:start
		
endclass:score_board


class environment;

        virtual inter.RM rm_inter;
        virtual inter.WM wm_inter;
        virtual inter.WD  wd_inter;	 

        mailbox #(packet) mgenwd = new;	
        mailbox #(packet) mwmrf  = new;
        mailbox #(packet) mrmsb  = new;
        mailbox #(packet) mrfsb  = new;
		
		function new(virtual inter.RM rm_inter,virtual inter.WM wm_inter,virtual inter.WD  wd_inter);
		              this.rm_inter = rm_inter;
					  this.wm_inter = wm_inter;
					  this.wd_inter = wd_inter;
		endfunction:new

        generator gen_h;
        write_drive wd_h;
        write_monitor wm_h;
        read_monitor rm_h;
        refence_model rf_h;
        score_board sb_h;
		
		
		
        task build();
              gen_h = new(mgenwd);
			  wd_h  = new(wd_inter,mgenwd);
			  wm_h  = new(wm_inter,mwmrf);
			  rm_h  = new(rm_inter,mrmsb);
              rf_h  = new(mwmrf,mrfsb);
              sb_h  = new(mrfsb,mrmsb);			  
        endtask:build	

       task start();
           gen_h.start();
           wd_h.start();
           wm_h.start();
           rm_h.start();
           rf_h.start();
           sb_h.start();
        endtask:start
		
		task stop();
		     wait(sb_h.DONE.triggered);
		endtask:stop	 

endclass:environment	

// classs test

class base_test;
    	 
        virtual inter.RM rm_inter;
        virtual inter.WM wm_inter;
        virtual inter.WD wd_inter;	
		
		environment env_h;
	    function new(virtual inter.RM rm_inter,virtual inter.WM wm_inter,virtual inter.WD wd_inter);
		              this.rm_inter = rm_inter;
					  this.wm_inter = wm_inter;
					  this.wd_inter = wd_inter;
					  env_h= new(rm_inter,wm_inter,wd_inter);
		endfunction:new
		 
        task build_and_start();

                env_h.build();
                env_h.start();
	        env_h.stop();
	        $finish;
        endtask:build_and_start   			 
  
endclass:base_test        

/*
class extend1 extends packet;

          constraint val_data1  { data_in inside{[2:5]};}


endclass:extend1

class base_extend1 extends base_test;

        

endclass:base_extend1

*/

module top;

      bit clk;
	  inter dut_if(clk);
	  
	  counter DUT(.clk(clk),.reset(dut_if.reset),.load(dut_if.load),.mode(dut_if.mode),.data_in(dut_if.data_in),.data_out(dut_if.data_out));

//module counter(clk,reset,load,mode,data_in,data_out);

	  
	  base_test bt;
	  
	  initial begin
	          bt = new (dut_if,dut_if,dut_if);
                  bt.build_and_start;
              end
           always #5 clk = ~clk;

endmodule:top 



/*

====================================== generator no_trans_id = 188======================================
                    0
no_load = 189 no_mode = 189 no_reset = 189

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 8 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 189======================================
                    0
no_load = 190 no_mode = 190 no_reset = 190

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 6 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 190======================================
                    0
no_load = 191 no_mode = 191 no_reset = 191

==================================== post randomize  t=0 ==================================================


 reset = 1 load = 0 data_in = 2 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 191======================================
                    0
no_load = 192 no_mode = 192 no_reset = 192

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 8 mode = 0


==============================================================================================================


====================================== generator no_trans_id = 192======================================
                    0
no_load = 193 no_mode = 193 no_reset = 193

==================================== post randomize  t=0 ==================================================


 reset = 1 load = 0 data_in = 9 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 193======================================
                    0
no_load = 194 no_mode = 194 no_reset = 194

==================================== post randomize  t=0 ==================================================


 reset = 1 load = 0 data_in = 5 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 194======================================
                    0
no_load = 195 no_mode = 195 no_reset = 195

==================================== post randomize  t=0 ==================================================


 reset = 1 load = 1 data_in = 0 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 195======================================
                    0
no_load = 196 no_mode = 196 no_reset = 196

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 0 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 196======================================
                    0
no_load = 197 no_mode = 197 no_reset = 197

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 0 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 197======================================
                    0
no_load = 198 no_mode = 198 no_reset = 198

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 0 data_in = 3 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 198======================================
                    0
no_load = 199 no_mode = 199 no_reset = 199

==================================== post randomize  t=0 ==================================================


 reset = 0 load = 1 data_in = 2 mode = 1


==============================================================================================================


====================================== generator no_trans_id = 199======================================
                    0
no_load = 200 no_mode = 200 no_reset = 200

==================================== post randomize  t=0 ==================================================


 reset = 1 load = 1 data_in = 10 mode = 0


==============================================================================================================


====================================== generator no_trans_id = 200======================================
                    0

====================================== Write Driver t=5 ======================================


====================================== Write Monitor t=5 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_in  = x

=========================================================================================================


====================================== Read Monitor t=5 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = x

=========================================================================================================


====================================== Refence Model t=5 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Compare is Failed
##########################################################################################

...............   30.000000  ................

====================================== Write Driver t=15 ======================================


====================================== Write Monitor t=15 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=15 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=15 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   43.571430  ................

====================================== Write Driver t=25 ======================================


====================================== Write Monitor t=25 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=25 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=25 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   53.571430  ................

====================================== Write Driver t=35 ======================================


====================================== Write Monitor t=35 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=35 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=35 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   53.571430  ................

====================================== Write Driver t=45 ======================================


====================================== Write Monitor t=45 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=45 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=45 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   53.571430  ................

====================================== Write Driver t=55 ======================================


====================================== Write Monitor t=55 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=55 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=55 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   64.285713  ................

====================================== Write Driver t=65 ======================================


====================================== Write Monitor t=65 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=65 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=65 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   64.285713  ................

====================================== Write Driver t=75 ======================================


====================================== Write Monitor t=75 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 11

=========================================================================================================


====================================== Read Monitor t=75 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=75 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   65.000000  ................

====================================== Write Driver t=85 ======================================


====================================== Write Monitor t=85 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=85 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=85 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   65.000000  ................

====================================== Write Driver t=95 ======================================


====================================== Write Monitor t=95 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=95 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 11

=========================================================================================================


====================================== Refence Model t=95 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 11

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   68.571426  ................

====================================== Write Driver t=105 ======================================


====================================== Write Monitor t=105 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_in  = 3

=========================================================================================================


====================================== Read Monitor t=105 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=105 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   69.285713  ................

====================================== Write Driver t=115 ======================================


====================================== Write Monitor t=115 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=115 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=115 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   69.285713  ................

====================================== Write Driver t=125 ======================================


====================================== Write Monitor t=125 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=125 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=125 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   69.285713  ................

====================================== Write Driver t=135 ======================================


====================================== Write Monitor t=135 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=135 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 2

=========================================================================================================


====================================== Refence Model t=135 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 2

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   72.857140  ................

====================================== Write Driver t=145 ======================================


====================================== Write Monitor t=145 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=145 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=145 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   72.857140  ................

====================================== Write Driver t=155 ======================================


====================================== Write Monitor t=155 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=155 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=155 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   72.857140  ................

====================================== Write Driver t=165 ======================================


====================================== Write Monitor t=165 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=165 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 2

=========================================================================================================


====================================== Refence Model t=165 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 2

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   73.571426  ................

====================================== Write Driver t=175 ======================================


====================================== Write Monitor t=175 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=175 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 3

=========================================================================================================


====================================== Refence Model t=175 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 3

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   74.285713  ................

====================================== Write Driver t=185 ======================================


====================================== Write Monitor t=185 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=185 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 8

=========================================================================================================


====================================== Refence Model t=185 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 8

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   81.428574  ................

====================================== Write Driver t=195 ======================================


====================================== Write Monitor t=195 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=195 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=195 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   81.428574  ................

====================================== Write Driver t=205 ======================================


====================================== Write Monitor t=205 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 11

=========================================================================================================


====================================== Read Monitor t=205 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=205 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   81.428574  ................

====================================== Write Driver t=215 ======================================


====================================== Write Monitor t=215 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=215 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


====================================== Refence Model t=215 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   82.142860  ................

====================================== Write Driver t=225 ======================================


====================================== Write Monitor t=225 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=225 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=225 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   82.142860  ................

====================================== Write Driver t=235 ======================================


====================================== Write Monitor t=235 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=235 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


====================================== Refence Model t=235 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   83.571426  ................

====================================== Write Driver t=245 ======================================


====================================== Write Monitor t=245 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=245 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=245 ======================================

 Reset = 0 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=255 ======================================


====================================== Write Monitor t=255 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_in  = 11

=========================================================================================================


====================================== Read Monitor t=255 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=255 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=265 ======================================


====================================== Write Monitor t=265 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 3

=========================================================================================================


====================================== Read Monitor t=265 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=265 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=275 ======================================


====================================== Write Monitor t=275 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=275 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=275 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=285 ======================================


====================================== Write Monitor t=285 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=285 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


====================================== Refence Model t=285 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=295 ======================================


====================================== Write Monitor t=295 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=295 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=295 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=305 ======================================


====================================== Write Monitor t=305 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=305 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=305 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=315 ======================================


====================================== Write Monitor t=315 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=315 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=315 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   84.285713  ................

====================================== Write Driver t=325 ======================================


====================================== Write Monitor t=325 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 3

=========================================================================================================


====================================== Read Monitor t=325 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 7

=========================================================================================================


====================================== Refence Model t=325 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 7

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=335 ======================================


====================================== Write Monitor t=335 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=335 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=335 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=345 ======================================


====================================== Write Monitor t=345 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=345 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=345 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=355 ======================================


====================================== Write Monitor t=355 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 4

=========================================================================================================


====================================== Read Monitor t=355 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


====================================== Refence Model t=355 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=365 ======================================


====================================== Write Monitor t=365 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 4

=========================================================================================================


====================================== Read Monitor t=365 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


====================================== Refence Model t=365 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=375 ======================================


====================================== Write Monitor t=375 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 4

=========================================================================================================


====================================== Read Monitor t=375 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=375 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=385 ======================================


====================================== Write Monitor t=385 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=385 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=385 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=395 ======================================


====================================== Write Monitor t=395 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=395 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=395 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=405 ======================================


====================================== Write Monitor t=405 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=405 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 2

=========================================================================================================


====================================== Refence Model t=405 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 2

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=415 ======================================


====================================== Write Monitor t=415 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=415 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 3

=========================================================================================================


====================================== Refence Model t=415 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 3

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   87.857147  ................

====================================== Write Driver t=425 ======================================


====================================== Write Monitor t=425 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=425 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 4

=========================================================================================================


====================================== Refence Model t=425 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 4

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=435 ======================================


====================================== Write Monitor t=435 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=435 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=435 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=445 ======================================


====================================== Write Monitor t=445 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 3

=========================================================================================================


====================================== Read Monitor t=445 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


====================================== Refence Model t=445 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=455 ======================================


====================================== Write Monitor t=455 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=455 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=455 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=465 ======================================


====================================== Write Monitor t=465 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=465 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=465 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=475 ======================================


====================================== Write Monitor t=475 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=475 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=475 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=485 ======================================


====================================== Write Monitor t=485 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=485 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=485 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=495 ======================================


====================================== Write Monitor t=495 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 4

=========================================================================================================


====================================== Read Monitor t=495 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=495 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=505 ======================================


====================================== Write Monitor t=505 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=505 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 4

=========================================================================================================


====================================== Refence Model t=505 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 4

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=515 ======================================


====================================== Write Monitor t=515 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=515 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 6

=========================================================================================================


====================================== Refence Model t=515 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 6

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   91.428574  ................

====================================== Write Driver t=525 ======================================


====================================== Write Monitor t=525 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=525 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 7

=========================================================================================================


====================================== Refence Model t=525 ======================================

 Reset = 0 Mode = 0  Load = 0 Data_out  = 7

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=535 ======================================


====================================== Write Monitor t=535 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=535 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=535 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=545 ======================================


====================================== Write Monitor t=545 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=545 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=545 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=555 ======================================


====================================== Write Monitor t=555 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=555 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=555 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=565 ======================================


====================================== Write Monitor t=565 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 4

=========================================================================================================


====================================== Read Monitor t=565 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=565 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=575 ======================================


====================================== Write Monitor t=575 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 5

=========================================================================================================


====================================== Read Monitor t=575 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


====================================== Refence Model t=575 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 11

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=585 ======================================


====================================== Write Monitor t=585 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=585 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=585 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=595 ======================================


====================================== Write Monitor t=595 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=595 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=595 ======================================

 Reset = 1 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=605 ======================================


====================================== Write Monitor t=605 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 6

=========================================================================================================


====================================== Read Monitor t=605 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=605 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=615 ======================================


====================================== Write Monitor t=615 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=615 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=615 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=625 ======================================


====================================== Write Monitor t=625 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 5

=========================================================================================================


====================================== Read Monitor t=625 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


====================================== Refence Model t=625 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 1

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   92.857140  ................

====================================== Write Driver t=635 ======================================


====================================== Write Monitor t=635 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=635 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 2

=========================================================================================================


====================================== Refence Model t=635 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 2

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=645 ======================================


====================================== Write Monitor t=645 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 10

=========================================================================================================


====================================== Read Monitor t=645 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=645 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=655 ======================================


====================================== Write Monitor t=655 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 7

=========================================================================================================


====================================== Read Monitor t=655 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


====================================== Refence Model t=655 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=665 ======================================


====================================== Write Monitor t=665 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=665 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=665 ======================================

 Reset = 0 Mode = 1  Load = 0 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=675 ======================================


====================================== Write Monitor t=675 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=675 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=675 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=685 ======================================


====================================== Write Monitor t=685 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 8

=========================================================================================================


====================================== Read Monitor t=685 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


====================================== Refence Model t=685 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 8

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=695 ======================================


====================================== Write Monitor t=695 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=695 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


====================================== Refence Model t=695 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=705 ======================================


====================================== Write Monitor t=705 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_in  = 1

=========================================================================================================


====================================== Read Monitor t=705 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=705 ======================================

 Reset = 1 Mode = 0  Load = 0 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=715 ======================================


====================================== Write Monitor t=715 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 0

=========================================================================================================


====================================== Read Monitor t=715 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


====================================== Refence Model t=715 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 9

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   93.571426  ................

====================================== Write Driver t=725 ======================================


====================================== Write Monitor t=725 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 3

=========================================================================================================


====================================== Read Monitor t=725 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 10

=========================================================================================================


====================================== Refence Model t=725 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 10

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   94.285713  ................

====================================== Write Driver t=735 ======================================


====================================== Write Monitor t=735 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_in  = 9

=========================================================================================================


====================================== Read Monitor t=735 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=735 ======================================

 Reset = 0 Mode = 1  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   94.285713  ................

====================================== Write Driver t=745 ======================================


====================================== Write Monitor t=745 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_in  = 5

=========================================================================================================


====================================== Read Monitor t=745 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


====================================== Refence Model t=745 ======================================

 Reset = 1 Mode = 0  Load = 1 Data_out  = 0

=========================================================================================================


##########################################################################################
                 Success Fully Compare
##########################################################################################

...............   94.285713  ................

====================================== Write Driver t=755 ======================================


====================================== Write Monitor t=755 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_in  = 2

=========================================================================================================


====================================== Read Monitor t=755 ======================================

 Reset = 1 Mode = 1  Load = 0 Data_out  = 5

==============================================================================

*/	  
       





      	   






					 
	  
      
	  

 			
         		  













 
         
