/********************************************************************************************

Copyright 2019 - Maven Silicon Softech Pvt Ltd.  
www.maven-silicon.com

All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.
It is not to be shared with or used by any third parties who have not enrolled for our paid 
training courses or received any written authorization from Maven Silicon.

Filename       :  ram_trans.sv   

Description    :  Transaction class for Dual Port Ram Testbench

Author Name    :  Putta Satish

Support e-mail :  techsupport_vm@maven-silicon.com 

Version        :  1.0

Date           :  02/06/2020

*********************************************************************************************/

// In class ram_trans

class ram_trans;     

   // Declare the following rand fields
     rand bit[64] data; 
   // data (bit/logic type , size 64)
     rand bit[12] rd_address,wr_address; 
   // rd_address, wr_address (bit/logic type , size 12)
     rand bit read,write; 
   // read, write (bit/logic type , size 1)     
     logic[64] data_out;
   // Declare a variable data_out (logic type , size 64)
        
   // Declare a static variable trans_id (int type), to keep the count of transactions generated
      static int trans_id;
        
   // Declare three static variables no_of_read_trans, no_of_write_trans, no_of_RW_trans (int type)
      static int  no_of_read_trans,no_of_write_trans,no_of_RW_trans; 

   // Add the following constraints 
   // wr_address!=rd_address;
 // read,write != 2'b00;

    constraint c {
                  wr_address != rd_address;  
                  {read,write} != 2'b00;  
                    data inside{[1:4294]}; 
                  } 
   // data between 1 and 4294   

     virtual function void display(input string a);
   //In virtual function display 
   // display the string         
   // display all the properties of the transaction class
     $display("\n####################################################################################################################################\n");
     $display("%s\t time = %t",a,$time);
     $display("write = %0d\twr_address = %0d\tdata = %0d\nread = %0d\trd_address = %0d\tdata_out = %0d",write,wr_address,data,read,rd_address,data_out); 
     $display("\n####################################################################################################################################\n");
     endfunction:display     

// In post_randomize method
      // Increment trans_id
      function void post_randomize;    
      // If it is only read transaction, increment no_of_read_trans
               if(this.read == 1'b1 && this.write == 1'b0)
                   no_of_read_trans++;       
      // If it is only write transaction, increment no_of_write_trans
               if(this.write == 1'b1 && this.read == 1'b0)
                   no_of_write_trans++;  
      // If it is read-write transaction, increment no_of_RW_trans
               if(this.read == 1'b1 && this.write == 1'b1)
                   no_of_RW_trans++;
      // call the display method and pass a string
              display("post_randomize ");
              $display("read trans = %0d , write trans = %0d , write and read = %0d ",no_of_read_trans,no_of_write_trans,no_of_RW_trans);  
       endfunction:post_randomize

endclass:ram_trans

/*
####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 1527	data = 2079
read = 1	rd_address = 3026	data_out = x

####################################################################################################################################

read trans = 1 , write trans = 0 , write and read = 0 

####################################################################################################################################

post_randomize 	 time =                41055
write = 1	wr_address = 2197	data = 3030
read = 0	rd_address = 28	data_out = x

####################################################################################################################################

read trans = 1 , write trans = 1 , write and read = 0 

####################################################################################################################################

post_randomize 	 time =                41055
write = 1	wr_address = 3650	data = 3843
read = 1	rd_address = 1017	data_out = x

####################################################################################################################################

read trans = 1 , write trans = 1 , write and read = 1 

####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 3088	data = 2801
read = 1	rd_address = 1901	data_out = x

####################################################################################################################################

read trans = 2 , write trans = 1 , write and read = 1 

####################################################################################################################################

post_randomize 	 time =                41055
write = 1	wr_address = 2926	data = 1841
read = 1	rd_address = 2038	data_out = x

####################################################################################################################################

read trans = 2 , write trans = 1 , write and read = 2 

####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 1366	data = 317
read = 1	rd_address = 1464	data_out = x

####################################################################################################################################

read trans = 3 , write trans = 1 , write and read = 2 

####################################################################################################################################

post_randomize 	 time =                41055
write = 1	wr_address = 3716	data = 1637
read = 1	rd_address = 1432	data_out = x

####################################################################################################################################

read trans = 3 , write trans = 1 , write and read = 3 

####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 2699	data = 3436
read = 1	rd_address = 2218	data_out = x

####################################################################################################################################

read trans = 4 , write trans = 1 , write and read = 3 

####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 554	data = 315
read = 1	rd_address = 1330	data_out = x

####################################################################################################################################

read trans = 5 , write trans = 1 , write and read = 3 

####################################################################################################################################

post_randomize 	 time =                41055
write = 0	wr_address = 1097	data = 1893
read = 1	rd_address = 2339	data_out = x

####################################################################################################################################

read trans = 6 , write trans = 1 , write and read = 3 

####################################################################################################################################

DATA FROM READ MONITOR	 time =                41075
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 3026	data_out = z

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41095
write = 0	wr_address = 0	data = 0
read = 0	rd_address = 3026	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41105
write = 1	wr_address = 2197	data = 3030
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41125
write = 0	wr_address = 2197	data = 3030
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41135
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 1017	data_out = z

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41145
write = 1	wr_address = 3650	data = 3843
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41155
write = 0	wr_address = 0	data = 0
read = 0	rd_address = 1017	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41175
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 1901	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41195
write = 1	wr_address = 2926	data = 1841
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41195
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 2038	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41215
write = 0	wr_address = 2926	data = 1841
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41215
write = 0	wr_address = 0	data = 0
read = 0	rd_address = 2038	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41235
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 1464	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41255
write = 1	wr_address = 3716	data = 1637
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41255
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 1432	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM WRITE MONITOR	 time =                41275
write = 0	wr_address = 3716	data = 1637
read = 0	rd_address = 0	data_out = x

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41275
write = 0	wr_address = 0	data = 0
read = 0	rd_address = 1432	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41295
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 2218	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41315
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 1330	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41335
write = 0	wr_address = 0	data = 0
read = 0	rd_address = 1330	data_out = 0

####################################################################################################################################


####################################################################################################################################

DATA FROM READ MONITOR	 time =                41355
write = 0	wr_address = 0	data = 0
read = 1	rd_address = 2339	data_out = 0

####################################################################################################################################

$finish called from file "../test/top.sv", line 70.
$finish at simulation time                42055
           V C S   S i m u l a t i o n   R e p o r t 
Time: 42055
*/
