





class trans;

        static  int i;
       static function  fun();
              int b;
               i++;
               b++;
          $display("\n*************************************************************************\n");
          $display(" value og b = %0d ,  i = %0d ", b,i);
          //$display("\n*************************************************************************\n");

        endfunction:fun
endclass:trans

  trans h,hb;
module test;

      initial begin
          // h = new;
          // hb =new;
           h.fun;
           h.fun;
           hb = h;
           hb.fun;
           //hb = new;
           //h = new;
           h.fun;
           hb.fun;
           h.fun;
           hb.fun;
        end
endmodule:test 


/*
output :
*************************************************************************

 value og b = 1 ,  i = 1 

*************************************************************************

 value og b = 1 ,  i = 2 

*************************************************************************

 value og b = 1 ,  i = 3 

*************************************************************************

 value og b = 1 ,  i = 4 

*************************************************************************

 value og b = 1 ,  i = 5 

*************************************************************************

 value og b = 1 ,  i = 6 

*************************************************************************

 value og b = 1 ,  i = 7 
           V C S   S i m u l a t i o n   R e p o r t 
*/
