


// creating  classes 

// grand parent class

class grandparent;
      virtual task send();
            $display("\n*******************************************************************************************\n");
            $display(" this is grand parent class ");
            $display("\n*******************************************************************************************\n");
      endtask:send
endclass:grandparent

// parent class 

class parent extends grandparent;
   
        virtual task send();
            $display("\n*******************************************************************************************\n");
            $display(" this is parent class ");
            $display("\n*******************************************************************************************\n");
        endtask:send

endclass:parent
                 
// child class

class child extends parent;
      
         virtual task send();
            $display("\n*******************************************************************************************\n");
            $display(" this is child  class ");
            $display("\n*******************************************************************************************\n");
          endtask:send
endclass:child  

// creating hanles fot child

   child ca,cb;
   parent pa,pb;
   grandparent ga,gb;

// creating the module for creating the object

module test;

      initial begin

           ca = new;
           //cb = new;
          
           pa = new;
           //pb = new;

           ga = new;
           //gb = new;

           ga.send;
           pa.send;
           ca.send;
           $display(" ****************** after pa = ca ****************************************************");
           pa = ca;
           pa.send; 
          $display(" ****************** after cb  = pa using $cast ****************************************");
            //cb = pa;
           $cast(cb,pa);         
           //cb = pa;
           cb.send;
           pa.send;
           pa = null;
           pa = new;
           pa.send;
           ga = pa;
           $display(" ****************** after ga = pa ****************************************************");
           ga.send;

           

       

        end

endmodule: test

 /*
*******************************************************************************************

 this is grand parent class 

*******************************************************************************************


*******************************************************************************************

 this is parent class 

*******************************************************************************************


*******************************************************************************************

 this is child  class 

*******************************************************************************************

 ****************** after pa = ca ****************************************************

*******************************************************************************************

 this is child  class 

*******************************************************************************************

 ****************** after cb  = pa using $cast ****************************************

*******************************************************************************************

 this is child  class 

*******************************************************************************************


*******************************************************************************************

 this is child  class 

*******************************************************************************************


*******************************************************************************************

 this is parent class 

*******************************************************************************************

 ****************** after ga = pa ****************************************************

*******************************************************************************************

 this is parent class 

*******************************************************************************************

           V C S   S i m u l a t i o n   R e p o r t 
*/    
 
