interface if3;
	logic a,b,c,d,e,f,i,j,k,l,m;
	modport moda(input a,d,e,f,h,output b,d,i,g);
	modport modb(input b,k,m,d,output c,j,a);
	modport modc(input g,h,
endinterface
