

// events checking 
// you have give lesser or equal vale where you used the @ or this wait then it triggered here we -> at #10 so you compulsary give lower then #10 for @ or //wait 

/*
module test;

    event ev;

      initial begin

           $display("\n########################################################################################################################\n");
           $display(" initial b1 drive control after 10 time units time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;

           $display("\n########################################################################################################################\n");
           $display(" initial b1 driving happening at time =%t ",$realtime);
           $display("\n########################################################################################################################\n");

           ->ev;
       end

      initial begin
           
           $display("\n########################################################################################################################\n");
           $display(" initial b2 about to drive  time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #9.4;
            //  #9.4 is consider as #9 and #9.5 abovr are consider as #10 

           @(ev);
           $display("\n########################################################################################################################\n");
           $display(" initial b2 data is driven at time =%t",$realtime);  
           $display("\n########################################################################################################################\n");

       end

endmodule:test       
*/
/*
if your givimng initial b2 as after #9 event triggerd 

########################################################################################################################

 initial b1 drive control after 10 time units time =                   0

########################################################################################################################


########################################################################################################################

 initial b2 about to drive  time =                   0

########################################################################################################################


########################################################################################################################

 initial b1 driving happening at time =                  10 

########################################################################################################################


########################################################################################################################

 initial b2 data is driven at time =                  10

########################################################################################################################

           V C S   S i m u l a t i o n   R e p o r t 

*/

/*
module test;

    event ev;

      initial begin

           $display("\n########################################################################################################################\n");
           $display(" initial b1 drive control after 10 time units time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;

           $display("\n########################################################################################################################\n");
           $display(" initial b1 driving happening at time =%t ",$realtime);
           $display("\n########################################################################################################################\n");

           ->ev;
       end

      initial begin
           
           $display("\n########################################################################################################################\n");
           $display(" initial b2 about to drive  time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;
            //  #9.4 is consider as #9 and #9.5 abovr are consider as #10 

           @(ev);
           $display("\n########################################################################################################################\n");
           $display(" initial b2 data is driven at time =%t",$realtime);  
           $display("\n########################################################################################################################\n");

       end

endmodule:test 

*/
/*

if your giving #10 for event this focus on  future  acope preset happend it cant be consderd so it is not display that
########################################################################################################################

 initial b1 drive control after 10 time units time =                   0

########################################################################################################################


########################################################################################################################

 initial b2 about to drive  time =                   0

########################################################################################################################


########################################################################################################################

 initial b1 driving happening at time =                  10 

########################################################################################################################

           V C S   S i m u l a t i o n   R e p o r t 
*/      

/*

module test;

    event ev;

      initial begin

           $display("\n########################################################################################################################\n");
           $display(" initial b1 drive control after 10 time units time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;

           $display("\n########################################################################################################################\n");
           $display(" initial b1 driving happening at time =%t ",$realtime);
           $display("\n########################################################################################################################\n");

           ->ev;
       end

      initial begin
           
           $display("\n########################################################################################################################\n");
           $display(" initial b2 about to drive  time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;
            //  #9.4 is consider as #9 and #9.5 abovr are consider as #10 

           wait(ev.triggered);
           $display("\n########################################################################################################################\n");
           $display(" initial b2 data is driven at time =%t",$realtime);  
           $display("\n########################################################################################################################\n");

       end

endmodule:test 

*/

/*

wait(ev.triggerd) is present and future scope so it consider both so its print 4 diplsays

########################################################################################################################

 initial b1 drive control after 10 time units time =                   0

########################################################################################################################


########################################################################################################################

 initial b2 about to drive  time =                   0

########################################################################################################################


########################################################################################################################

 initial b1 driving happening at time =                  10 

########################################################################################################################


########################################################################################################################

 initial b2 data is driven at time =                  10

########################################################################################################################

           V C S   S i m u l a t i o n   R e p o r t 

*/

module test;

    event ev;

      initial begin

           $display("\n########################################################################################################################\n");
           $display(" initial b1 drive control after 10 time units time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10;

           $display("\n########################################################################################################################\n");
           $display(" initial b1 driving happening at time =%t ",$realtime);
           $display("\n########################################################################################################################\n");

           ->ev;
       end

      initial begin
           
           $display("\n########################################################################################################################\n");
           $display(" initial b2 about to drive  time =%t",$realtime);
           $display("\n########################################################################################################################\n");

           #10.3;
            //  #9.4 is consider as #9 and #9.5 abovr are consider as #10 

           wait(ev.triggered);
           $display("\n########################################################################################################################\n");
           $display(" initial b2 data is driven at time =%t",$realtime);  
           $display("\n########################################################################################################################\n");

       end

endmodule:test 

/*
########################################################################################################################

 initial b1 drive control after 10 time units time =                   0

########################################################################################################################


########################################################################################################################

 initial b2 about to drive  time =                   0

########################################################################################################################


########################################################################################################################

 initial b1 driving happening at time =                  10 

########################################################################################################################


########################################################################################################################

 initial b2 data is driven at time =                  10

########################################################################################################################

           V C S   S i m u l a t i o n   R e p o r t 
*/


