

module arrays();

// declaring the packed arrays 

     bit [7:0][3:0] packed_nibble; // 8 nibbles into 32 bit
// first vector gives you number of groups and second vector gives number of bits per each group 

     bit [3:0][7:0] packed_byte; // 4 bytes into 32 bits 4*8=32
  
     initial
            begin
                 $display("============================================================================================================================");
                 packed_nibble = 32'hABCD_1234;
                 packed_byte = 32'hABCD_1234;
                 $display("total_packet nibble = %b \n, least significant nibble =%b \n,0'rth lsb  bit of least signficant nibble=%b "
,packed_nibble,packed_nibble[7],packed_nibble[7][0]);
                 $display("total_packet byte = %b \n , least significant byte =%b \n,0'rth lsb bit of least signficant byte=%b "
,packed_byte,packed_byte[3],packed_byte[3][0]);
          $display("============================================================================================================================");


            end

// declaring the unpacked array of 3 packed elemnts

  bit [3:0] [7:0] bytes [0:2];
  

  initial begin
       
      #30;
        $display("============================================================================================================================");

      bytes[0]=32'd255;
       $display(" totoal packet = %p ",bytes);
        $display(" totoal 0 rth element = %b ",bytes[0]);

      // assinging the 0 rth element
     bytes[0][3] = 32'd20;
      $display(" 0 rth element and 3rd group = %b ",bytes[0][3]);
      // asssiging the 0 rth element and 3rd group byte
     bytes[0][3][6]=1'b0; 
      $display(" orth element 3rd group 6th bit = %b ", bytes[0][3][6]);          
      // assinging the 0 rth element  and 3rd gruop and 6th bit 
     $display("============================================================================================================================");

      end
   
// accesssing the elements of array

     int  mdst[3][5] = '{'{01,21,32,34,45},'{123,323,43,54,34},'{123,345,64,57,67}};
      
 
     initial begin
      #60;
    $display("============================================================================================================================");

     // for (int i=0;i<$size(msrc);i++)
         //  msrc[i]=i;
     $display(" totoal  = %p ",mdst);

      foreach(mdst[i,j])
          $display("mdst[%0d][%0d] = %0d",i,j,mdst[i][j]); 
     $display("============================================================================================================================");
   
     end    
//  aggregate  copy & compare

     bit [31:0] ms[5] = '{0,1,2,3,4},mt[5] = '{5,4,3,2,1};
    initial begin
    #80;
   $display("============================================================================================================================");

     if(ms == mt)
       $display(" ms=%p is equal to mt=%p ",ms,mt);
     else
       $display(" ms=%p is not equal to mt=p ",ms,mt);

    ms =mt;

    if(ms [1:4] == mt[1:4])  
       $display(" ms[1:4]=%p is equal to mt[1:4]=%p ",ms[1:4],mt[1:4]);
    else
       $display(" ms[1:4]=%p is not equal to mt[1:4]=%p ",ms[1:4],mt[1:4]);
   $display("============================================================================================================================");

    end

// dynamic array 

   int da1[],da2[];

     initial begin
     #100
     $display("============================================================================================================================");
     da1 = new[20];
     foreach(da1[i])
        da1[i]=i;
     $display(" da1[10]=%p ",da1); 
     da2=da1;
     da1 =new[30](da1);
         $display(" da1[30]=%p ",da1); 
    $display(" da2[10]=%p ",da2); 
     da2.delete();
      $display("da2 = %p ",da2);
       $display(" da1[30]=%p ",da1);
     $display("============================================================================================================================");
     end 

// queues  

   int qm1[$] = '{1,3,4,5,6};
   int qm2[$] =  '{2,3};
   int k = 32;
   initial begin
   #120;
   $display("============================================================================================================================");
    
   qm1.insert(1,k);
   qm1.delete(1);
   qm1.push_back(40);
   qm1.push_front(8);
   $display("qm1 = %p " ,qm1);
   $display("qm2 = %p " ,qm2);
   k=qm1.pop_back();
    $display("qm1 = %p " ,qm1);

    qm2.push_back(12);
 $display("qm2 = %p " ,qm2);

   k=qm2.pop_front(); 
   $display("qm2 = %p " ,qm2);
   foreach(qm1[i])
    $display(qm1[i]);
    qm2.delete();
   $display("============================================================================================================================");
   end  
   
endmodule      


/*

OUTPUT :

============================================================================================================================
# total_packet nibble = 10101011110011010001001000110100 
# , least significant nibble =1010 
# ,0'rth lsb  bit of least signficant nibble=0 
# total_packet byte = 10101011110011010001001000110100 
#  , least significant byte =10101011 
# ,0'rth lsb bit of least signficant byte=1 
# ============================================================================================================================
# ============================================================================================================================
#  totoal packet = '{'{0, 0, 0, 255}, '{0, 0, 0, 0}, '{0, 0, 0, 0}} 
#  totoal 0 rth element = 00000000000000000000000011111111 
#  0 rth element and 3rd group = 00010100 
#  orth element 3rd group 6th bit = 0 
# ============================================================================================================================
# ============================================================================================================================
#  totoal  = '{'{1, 21, 32, 34, 45}, '{123, 323, 43, 54, 34}, '{123, 345, 64, 57, 67}} 
# mdst[0][0] = 1
# mdst[0][1] = 21
# mdst[0][2] = 32
# mdst[0][3] = 34
# mdst[0][4] = 45
# mdst[1][0] = 123
# mdst[1][1] = 323
# mdst[1][2] = 43
# mdst[1][3] = 54
# mdst[1][4] = 34
# mdst[2][0] = 123
# mdst[2][1] = 345
# mdst[2][2] = 64
# mdst[2][3] = 57
# mdst[2][4] = 67
# ============================================================================================================================
# ============================================================================================================================
#  ms='{0, 1, 2, 3, 4} is not equal to mt=p 
#  ms[1:4]='{4, 3, 2, 1} is equal to mt[1:4]='{4, 3, 2, 1} 
# ============================================================================================================================
# ============================================================================================================================
#  da1[10]='{0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19} 
#  da1[30]='{0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0} 
#  da2[10]='{0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19} 
# da2 = '{} 
#  da1[30]='{0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0} 
# ============================================================================================================================
# ============================================================================================================================
# qm1 = '{8, 1, 3, 4, 5, 6, 40} 
# qm2 = '{2, 3} 
# qm1 = '{8, 1, 3, 4, 5, 6} 
# qm2 = '{2, 3, 12} 
# qm2 = '{3, 12} 
#           8
#           1
#           3
#           4
#           5
#           6
# ============================================================================================================================

*/  
