

module test_semaphore;

	// In class driver
 
class driver;
            
		// write task send with input argument of string type
      task send(input string a);
             
			// Get the key using sem handle 

             sem.get(1);

			// Display the string which indicates the respective driver information
             $display("\n*******************************************************************************************\n");
             $display(" time = %0t -- put -- handle = %s",$time,a);
             $display("\n*******************************************************************************************\n");
             #10;
 
			// Put the key using sem handle 

           // sem.put(1);

			// Display the string which indicates the respective driver information
             $display(" \n*******************************************************************************************\n");
             $display(" time = %0t -- get -- handle = %s",$time,a);
             $display("\n*******************************************************************************************\n");

        endtask:send 
endclass:driver

	// Declare an array of two drivers  
          
driver da[2];

semaphore sem;
    
           
	// Declare a handle for semaphore

	// Within initial block
               initial begin
		// Create instances of drivers
                 da[0]  =  new;
                 da[1]  =  new;

		// Create the instance of semaphore handle and initialize it with 1 key
                sem = new(0);


		// Call send task of both drivers 5 times within fork join
                fork 
                da[0].send("da[0]");
                da[0].send("da[0]");
                da[1].send("da[1]");
                da[1].send("da[1]");
                da[0].send("da[0]");
                da[1].send("da[1]");


                join
		// pass any meaning full string message to indicate the driver information
                $display("\n*******************************************************************************************\n");
                $display("\nda[0] = %0p\nda[1] = %0p\n",da[0],da[1]);
                $display("\n*******************************************************************************************\n");

                end
	endmodule 


/*

// yout giving only kew token but here you called 5 threads inside so first thread get key and wait put the key token 
// if get key tokens will decremented like this ways if you put key token incresed 

//  sem = new(1);
//  sem.get(1);
//  sem.put(1);


*******************************************************************************************

 time = 0 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 20 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 20 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 30 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 30 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 40 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 40 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 50 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 50 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 60 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************


da[0] = '{}
da[1] = '{}


*******************************************************************************************

           V C S   S i m u l a t i o n   R e p o r t 

*/


/*

//when i was not givng put and gving 

// all are excute normal forkjoin  #0 first diplay of get  first 3 and #10 display of put first 3
                da[0].send("da[0]");
                da[0].send("da[0]");
                da[1].send("da[1]");
// these will excuted it takes the 3 key tokens 

// if your calling 3 threads inside a fork join you giving 3 tokens in sem = new (3) they not waiting for putting sufficent token are there so all are excu//ted parallel 

// sem = new(3);

//sem.get(1);


                fork 
                da[0].send("da[0]");
                da[0].send("da[0]");
                da[1].send("da[1]");

                da[1].send("da[1]");
                da[0].send("da[0]");
                da[1].send("da[1]");
                join

*******************************************************************************************

 time = 0 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- put -- handle = da[1]

*******************************************************************************************

           V C S   S i m u l a t i o n   R e p o r t 


*/

/*

//when i was not givng put and gving 

// sem = new(3);

//sem.get(3);
                fork 
                da[0].send("da[0]");

                da[0].send("da[0]");
                da[1].send("da[1]");
                da[1].send("da[1]");
                da[0].send("da[0]");
                da[1].send("da[1]");
                join


*******************************************************************************************

 time = 0 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- put -- handle = da[0]

*******************************************************************************************

           V C S   S i m u l a t i o n   R e p o r t 
*/


/*

//if your giving put key token first then get key token 

// all the threads working parallel beacuse each thred going task same time but due to number of key tokens they waited but here you givng put(1)
// each thered givnig their own thread so all are accesing same time  


 sem.put(1);

 sem.get(1);

 sem = new(0);

                fork 
                da[0].send("da[0]");
                da[0].send("da[0]");
                da[1].send("da[1]");
                da[1].send("da[1]");
                da[0].send("da[0]");
                da[1].send("da[1]");
                join

*******************************************************************************************

 time = 0 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- put -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 0 -- put -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[0]

*******************************************************************************************


*******************************************************************************************

 time = 10 -- get -- handle = da[1]

*******************************************************************************************


*******************************************************************************************


da[0] = '{}
da[1] = '{}


*******************************************************************************************

           V C S   S i m u l a t i o n   R e p o r t 

*/






